Transfer Function Analysis
*By Chris Vasquez

.lib "nom.lib" 

*Analysis directives: 
.TF V([2]) V_V2
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 



**** INCLUDING SCHEMATIC1.net ****
* source VOLTAGE AMPLIFIER
.EXTERNAL OUTPUT 2
.EXTERNAL OUTPUT 1
Q_Q4         2 1 N47435 Q2N2222
R_R3         0 1 R_R3 100k TC=25PPM,0 
.model        R_R3 RES R=1 DEV=0.1% TC1=25PPM TC2=0
R_R4         0 N47435 R_R4 400 TC=25PPM,0 
.model        R_R4 RES R=1 DEV=0.1% TC1=25PPM TC2=0
R_R2         2 N47261 R_R2 3k TC=50PPM,0 
.model        R_R2 RES R=1 DEV=0.1% TC1=50PPM TC2=0
C_C2         0 N47435  330u  TC=0,0 
R_R1         1 N47261 R_R1 300k TC=25PPM,0 
.model        R_R1 RES R=1 DEV=0.1% TC1=25PPM TC2=0
V_V1         N47407 0  AC 0.01
+SIN 0 0 1k 0 0 0
C_C1         1 N47407  330u  TC=0,0 
V_V2         N47261 0 9Vdc

**** RESUMING sim.cir ****
.END

**** 04/30/20 15:34:14 ****** PSpice 17.2.0 (March 2016) ****** ID# 0 ********

 ** Profile: "SCHEMATIC1-sim"  [ c:\users\chris\documents\pspice\voltage amplifier-pspicefiles\schematic1\sim.sim ] 


 ****     BJT MODEL PARAMETERS


******************************************************************************




               Q2N2222         
               NPN             
       LEVEL    1            
          IS   14.340000E-15 
          BF  255.9          
          NF    1            
         VAF   74.03         
         IKF     .2847       
         ISE   14.340000E-15 
          NE    1.307        
          BR    6.092        
          NR    1            
         ISS    0            
          RB   10            
          RE    0            
          RC    1            
         CJE   22.010000E-12 
         VJE     .75         
         MJE     .377        
         CJC    7.306000E-12 
         VJC     .75         
         MJC     .3416       
        XCJC    1            
         CJS    0            
         VJS     .75         
          TF  411.100000E-12 
         XTF    3            
         VTF    1.7          
         ITF     .6          
          TR   46.910000E-09 
         XTB    1.5          
          KF    0            
          AF    1            
          CN    2.42         
           D     .87         


**** 04/30/20 15:34:14 ****** PSpice 17.2.0 (March 2016) ****** ID# 0 ********

 ** Profile: "SCHEMATIC1-sim"  [ c:\users\chris\documents\pspice\voltage amplifier-pspicefiles\schematic1\sim.sim ] 


 ****     Resistor MODEL PARAMETERS


******************************************************************************




               R_R3            R_R4            R_R2            R_R1            
           R    1               1               1               1            
         TC1   25.000000E-12   25.000000E-12   50.000000E-12   25.000000E-12 


**** 04/30/20 15:34:14 ****** PSpice 17.2.0 (March 2016) ****** ID# 0 ********

 ** Profile: "SCHEMATIC1-sim"  [ c:\users\chris\documents\pspice\voltage amplifier-pspicefiles\schematic1\sim.sim ] 


 ****     SMALL SIGNAL BIAS SOLUTION       TEMPERATURE =   27.000 DEG C


******************************************************************************



 NODE   VOLTAGE     NODE   VOLTAGE     NODE   VOLTAGE     NODE   VOLTAGE


(    1)    1.3953  (    2)    3.5257  (N47261)    9.0000 (N47407)    0.0000     

(N47435)     .7345 




    VOLTAGE SOURCE CURRENTS
    NAME         CURRENT

    V_V1         0.000E+00
    V_V2        -1.850E-03

    TOTAL POWER DISSIPATION   1.67E-02  WATTS






 ****     SMALL-SIGNAL CHARACTERISTICS


      V(2)/V_V2 =  1.128E-01

      INPUT RESISTANCE AT V_V2 =  3.348E+03

      OUTPUT RESISTANCE AT V(2) =  2.891E+03


          JOB CONCLUDED

**** 04/30/20 15:34:14 ****** PSpice 17.2.0 (March 2016) ****** ID# 0 ********

 ** Profile: "SCHEMATIC1-sim"  [ c:\users\chris\documents\pspice\voltage amplifier-pspicefiles\schematic1\sim.sim ] 


 ****     JOB STATISTICS SUMMARY


******************************************************************************



  License check-out time            =        1.45
  Total job time (using Solver 1)   =         .05
